module HPC2(
    clk,
    a0,
    a1,
    a2,
    a3,
    a4,
    b0,
    b1,
    b2,
    b3,
    b4,
    r01,
    r02,
    r03,
    r04,
    r12,
    r13,
    r14,
    r23,
    r24,
    r34,
    c0,
    c1,
    c2,
    c3,
    c4,
);
//INPUTS
    input clk;
    input  [7:0] a0;
    input  [7:0] a1;
    input  [7:0] a2;
    input  [7:0] a3;
    input  [7:0] a4;
    input  [7:0] b0;
    input  [7:0] b1;
    input  [7:0] b2;
    input  [7:0] b3;
    input  [7:0] b4;
    input  [7:0] r01;
    input  [7:0] r02;
    input  [7:0] r03;
    input  [7:0] r04;
    input  [7:0] r12;
    input  [7:0] r13;
    input  [7:0] r14;
    input  [7:0] r23;
    input  [7:0] r24;
    input  [7:0] r34;
//OUTPUTS
    output reg  [7:0] c0;
    output reg  [7:0] c1;
    output reg  [7:0] c2;
    output reg  [7:0] c3;
    output reg  [7:0] c4;
//Intermediate values
    wire [7:0] a0_inp;
    wire [7:0] a1_inp;
    wire [7:0] a2_inp;
    wire [7:0] a3_inp;
    wire [7:0] a4_inp;
    wire [7:0] b0_inp;
    wire [7:0] b1_inp;
    wire [7:0] b2_inp;
    wire [7:0] b3_inp;
    wire [7:0] b4_inp;
    wire [7:0] r01_inp;
    wire [7:0] r02_inp;
    wire [7:0] r03_inp;
    wire [7:0] r04_inp;
    wire [7:0] r12_inp;
    wire [7:0] r13_inp;
    wire [7:0] r14_inp;
    wire [7:0] r23_inp;
    wire [7:0] r24_inp;
    wire [7:0] r34_inp;
    reg [7:0] b_share_reg_hpc2_same_shares_4_order0;
    reg [7:0] a0_inp_reg;
    wire [7:0] z1_assgn1;
    reg [7:0] u00;
    reg [7:0] temp_hpc2_v_4_order0;
    wire [7:0] z3_assgn3;
    reg [7:0] v01;
    reg [7:0] rand_reg_hpc2_w_4_order0;
    wire [7:0] a_neg_hpc2_w_4_order0;
    reg [7:0] a_neg_hpc2_w_4_order0_reg;
    wire [7:0] z5_assgn5;
    reg [7:0] w01;
    wire [7:0] u01;
    reg [7:0] temp_hpc2_v_4_order1;
    wire [7:0] z7_assgn7;
    reg [7:0] v02;
    reg [7:0] rand_reg_hpc2_w_4_order1;
    wire [7:0] a_neg_hpc2_w_4_order1;
    reg [7:0] a_neg_hpc2_w_4_order1_reg;
    wire [7:0] z9_assgn9;
    reg [7:0] w02;
    wire [7:0] u02;
    reg [7:0] temp_hpc2_v_4_order2;
    wire [7:0] z11_assgn11;
    reg [7:0] v03;
    reg [7:0] rand_reg_hpc2_w_4_order2;
    wire [7:0] a_neg_hpc2_w_4_order2;
    reg [7:0] a_neg_hpc2_w_4_order2_reg;
    wire [7:0] z13_assgn13;
    reg [7:0] w03;
    wire [7:0] u03;
    reg [7:0] temp_hpc2_v_4_order3;
    wire [7:0] z15_assgn15;
    reg [7:0] v04;
    reg [7:0] rand_reg_hpc2_w_4_order3;
    wire [7:0] a_neg_hpc2_w_4_order3;
    reg [7:0] a_neg_hpc2_w_4_order3_reg;
    wire [7:0] z17_assgn17;
    reg [7:0] w04;
    wire [7:0] u04;
    reg [7:0] temp_hpc2_v_4_order4;
    reg [7:0] a1_inp_reg;
    wire [7:0] z19_assgn19;
    reg [7:0] v10;
    reg [7:0] rand_reg_hpc2_w_4_order4;
    wire [7:0] a_neg_hpc2_w_4_order4;
    reg [7:0] a_neg_hpc2_w_4_order4_reg;
    wire [7:0] z21_assgn21;
    reg [7:0] w10;
    wire [7:0] u10;
    reg [7:0] b_share_reg_hpc2_same_shares_4_order1;
    wire [7:0] z23_assgn23;
    reg [7:0] u11;
    reg [7:0] temp_hpc2_v_4_order5;
    wire [7:0] z25_assgn25;
    reg [7:0] v12;
    reg [7:0] rand_reg_hpc2_w_4_order5;
    wire [7:0] a_neg_hpc2_w_4_order5;
    reg [7:0] a_neg_hpc2_w_4_order5_reg;
    wire [7:0] z27_assgn27;
    reg [7:0] w12;
    wire [7:0] u12;
    reg [7:0] temp_hpc2_v_4_order6;
    wire [7:0] z29_assgn29;
    reg [7:0] v13;
    reg [7:0] rand_reg_hpc2_w_4_order6;
    wire [7:0] a_neg_hpc2_w_4_order6;
    reg [7:0] a_neg_hpc2_w_4_order6_reg;
    wire [7:0] z31_assgn31;
    reg [7:0] w13;
    wire [7:0] u13;
    reg [7:0] temp_hpc2_v_4_order7;
    wire [7:0] z33_assgn33;
    reg [7:0] v14;
    reg [7:0] rand_reg_hpc2_w_4_order7;
    wire [7:0] a_neg_hpc2_w_4_order7;
    reg [7:0] a_neg_hpc2_w_4_order7_reg;
    wire [7:0] z35_assgn35;
    reg [7:0] w14;
    wire [7:0] u14;
    reg [7:0] temp_hpc2_v_4_order8;
    reg [7:0] a2_inp_reg;
    wire [7:0] z37_assgn37;
    reg [7:0] v20;
    reg [7:0] rand_reg_hpc2_w_4_order8;
    wire [7:0] a_neg_hpc2_w_4_order8;
    reg [7:0] a_neg_hpc2_w_4_order8_reg;
    wire [7:0] z39_assgn39;
    reg [7:0] w20;
    wire [7:0] u20;
    reg [7:0] temp_hpc2_v_4_order9;
    wire [7:0] z41_assgn41;
    reg [7:0] v21;
    reg [7:0] rand_reg_hpc2_w_4_order9;
    wire [7:0] a_neg_hpc2_w_4_order9;
    reg [7:0] a_neg_hpc2_w_4_order9_reg;
    wire [7:0] z43_assgn43;
    reg [7:0] w21;
    wire [7:0] u21;
    reg [7:0] b_share_reg_hpc2_same_shares_4_order2;
    wire [7:0] z45_assgn45;
    reg [7:0] u22;
    reg [7:0] temp_hpc2_v_4_order10;
    wire [7:0] z47_assgn47;
    reg [7:0] v23;
    reg [7:0] rand_reg_hpc2_w_4_order10;
    wire [7:0] a_neg_hpc2_w_4_order10;
    reg [7:0] a_neg_hpc2_w_4_order10_reg;
    wire [7:0] z49_assgn49;
    reg [7:0] w23;
    wire [7:0] u23;
    reg [7:0] temp_hpc2_v_4_order11;
    wire [7:0] z51_assgn51;
    reg [7:0] v24;
    reg [7:0] rand_reg_hpc2_w_4_order11;
    wire [7:0] a_neg_hpc2_w_4_order11;
    reg [7:0] a_neg_hpc2_w_4_order11_reg;
    wire [7:0] z53_assgn53;
    reg [7:0] w24;
    wire [7:0] u24;
    reg [7:0] temp_hpc2_v_4_order12;
    reg [7:0] a3_inp_reg;
    wire [7:0] z55_assgn55;
    reg [7:0] v30;
    reg [7:0] rand_reg_hpc2_w_4_order12;
    wire [7:0] a_neg_hpc2_w_4_order12;
    reg [7:0] a_neg_hpc2_w_4_order12_reg;
    wire [7:0] z57_assgn57;
    reg [7:0] w30;
    wire [7:0] u30;
    reg [7:0] temp_hpc2_v_4_order13;
    wire [7:0] z59_assgn59;
    reg [7:0] v31;
    reg [7:0] rand_reg_hpc2_w_4_order13;
    wire [7:0] a_neg_hpc2_w_4_order13;
    reg [7:0] a_neg_hpc2_w_4_order13_reg;
    wire [7:0] z61_assgn61;
    reg [7:0] w31;
    wire [7:0] u31;
    reg [7:0] temp_hpc2_v_4_order14;
    wire [7:0] z63_assgn63;
    reg [7:0] v32;
    reg [7:0] rand_reg_hpc2_w_4_order14;
    wire [7:0] a_neg_hpc2_w_4_order14;
    reg [7:0] a_neg_hpc2_w_4_order14_reg;
    wire [7:0] z65_assgn65;
    reg [7:0] w32;
    wire [7:0] u32;
    reg [7:0] b_share_reg_hpc2_same_shares_4_order3;
    wire [7:0] z67_assgn67;
    reg [7:0] u33;
    reg [7:0] temp_hpc2_v_4_order15;
    wire [7:0] z69_assgn69;
    reg [7:0] v34;
    reg [7:0] rand_reg_hpc2_w_4_order15;
    wire [7:0] a_neg_hpc2_w_4_order15;
    reg [7:0] a_neg_hpc2_w_4_order15_reg;
    wire [7:0] z71_assgn71;
    reg [7:0] w34;
    wire [7:0] u34;
    reg [7:0] temp_hpc2_v_4_order16;
    reg [7:0] a4_inp_reg;
    wire [7:0] z73_assgn73;
    reg [7:0] v40;
    reg [7:0] rand_reg_hpc2_w_4_order16;
    wire [7:0] a_neg_hpc2_w_4_order16;
    reg [7:0] a_neg_hpc2_w_4_order16_reg;
    wire [7:0] z75_assgn75;
    reg [7:0] w40;
    wire [7:0] u40;
    reg [7:0] temp_hpc2_v_4_order17;
    wire [7:0] z77_assgn77;
    reg [7:0] v41;
    reg [7:0] rand_reg_hpc2_w_4_order17;
    wire [7:0] a_neg_hpc2_w_4_order17;
    reg [7:0] a_neg_hpc2_w_4_order17_reg;
    wire [7:0] z79_assgn79;
    reg [7:0] w41;
    wire [7:0] u41;
    reg [7:0] temp_hpc2_v_4_order18;
    wire [7:0] z81_assgn81;
    reg [7:0] v42;
    reg [7:0] rand_reg_hpc2_w_4_order18;
    wire [7:0] a_neg_hpc2_w_4_order18;
    reg [7:0] a_neg_hpc2_w_4_order18_reg;
    wire [7:0] z83_assgn83;
    reg [7:0] w42;
    wire [7:0] u42;
    reg [7:0] temp_hpc2_v_4_order19;
    wire [7:0] z85_assgn85;
    reg [7:0] v43;
    reg [7:0] rand_reg_hpc2_w_4_order19;
    wire [7:0] a_neg_hpc2_w_4_order19;
    reg [7:0] a_neg_hpc2_w_4_order19_reg;
    wire [7:0] z87_assgn87;
    reg [7:0] w43;
    wire [7:0] u43;
    reg [7:0] b_share_reg_hpc2_same_shares_4_order4;
    wire [7:0] z89_assgn89;
    reg [7:0] u44;
    wire [7:0] t1;
    wire [7:0] t2;
    wire [7:0] t3;
    wire [7:0] t4;
    wire [7:0] t5;
    wire [7:0] t6;
    wire [7:0] t7;
    wire [7:0] t8;
    wire [7:0] t9;
    wire [7:0] t10;
    wire [7:0] t11;
    wire [7:0] t12;
    wire [7:0] t13;
    wire [7:0] t14;
    wire [7:0] t15;

    assign a0_inp = a0;
    assign a1_inp = a1;
    assign a2_inp = a2;
    assign a3_inp = a3;
    assign a4_inp = a4;
    assign b0_inp = b0;
    assign b1_inp = b1;
    assign b2_inp = b2;
    assign b3_inp = b3;
    assign b4_inp = b4;
    assign r01_inp = r01;
    assign r02_inp = r02;
    assign r03_inp = r03;
    assign r04_inp = r04;
    assign r12_inp = r12;
    assign r13_inp = r13;
    assign r14_inp = r14;
    assign r23_inp = r23;
    assign r24_inp = r24;
    assign r34_inp = r34;
    assign z1_assgn1 = (a0_inp_reg & b_share_reg_hpc2_same_shares_4_order0);
    assign z3_assgn3 = (temp_hpc2_v_4_order0 & a0_inp_reg);
    assign a_neg_hpc2_w_4_order0 = !a0_inp;
    assign z5_assgn5 = (a_neg_hpc2_w_4_order0_reg & rand_reg_hpc2_w_4_order0);
    assign u01 = (v01 ^ w01);
    assign z7_assgn7 = (temp_hpc2_v_4_order1 & a0_inp_reg);
    assign a_neg_hpc2_w_4_order1 = !a0_inp;
    assign z9_assgn9 = (a_neg_hpc2_w_4_order1_reg & rand_reg_hpc2_w_4_order1);
    assign u02 = (v02 ^ w02);
    assign z11_assgn11 = (temp_hpc2_v_4_order2 & a0_inp_reg);
    assign a_neg_hpc2_w_4_order2 = !a0_inp;
    assign z13_assgn13 = (a_neg_hpc2_w_4_order2_reg & rand_reg_hpc2_w_4_order2);
    assign u03 = (v03 ^ w03);
    assign z15_assgn15 = (temp_hpc2_v_4_order3 & a0_inp_reg);
    assign a_neg_hpc2_w_4_order3 = !a0_inp;
    assign z17_assgn17 = (a_neg_hpc2_w_4_order3_reg & rand_reg_hpc2_w_4_order3);
    assign u04 = (v04 ^ w04);
    assign z19_assgn19 = (temp_hpc2_v_4_order4 & a1_inp_reg);
    assign a_neg_hpc2_w_4_order4 = !a1_inp;
    assign z21_assgn21 = (a_neg_hpc2_w_4_order4_reg & rand_reg_hpc2_w_4_order4);
    assign u10 = (v10 ^ w10);
    assign z23_assgn23 = (a1_inp_reg & b_share_reg_hpc2_same_shares_4_order1);
    assign z25_assgn25 = (temp_hpc2_v_4_order5 & a1_inp_reg);
    assign a_neg_hpc2_w_4_order5 = !a1_inp;
    assign z27_assgn27 = (a_neg_hpc2_w_4_order5_reg & rand_reg_hpc2_w_4_order5);
    assign u12 = (v12 ^ w12);
    assign z29_assgn29 = (temp_hpc2_v_4_order6 & a1_inp_reg);
    assign a_neg_hpc2_w_4_order6 = !a1_inp;
    assign z31_assgn31 = (a_neg_hpc2_w_4_order6_reg & rand_reg_hpc2_w_4_order6);
    assign u13 = (v13 ^ w13);
    assign z33_assgn33 = (temp_hpc2_v_4_order7 & a1_inp_reg);
    assign a_neg_hpc2_w_4_order7 = !a1_inp;
    assign z35_assgn35 = (a_neg_hpc2_w_4_order7_reg & rand_reg_hpc2_w_4_order7);
    assign u14 = (v14 ^ w14);
    assign z37_assgn37 = (temp_hpc2_v_4_order8 & a2_inp_reg);
    assign a_neg_hpc2_w_4_order8 = !a2_inp;
    assign z39_assgn39 = (a_neg_hpc2_w_4_order8_reg & rand_reg_hpc2_w_4_order8);
    assign u20 = (v20 ^ w20);
    assign z41_assgn41 = (temp_hpc2_v_4_order9 & a2_inp_reg);
    assign a_neg_hpc2_w_4_order9 = !a2_inp;
    assign z43_assgn43 = (a_neg_hpc2_w_4_order9_reg & rand_reg_hpc2_w_4_order9);
    assign u21 = (v21 ^ w21);
    assign z45_assgn45 = (a2_inp_reg & b_share_reg_hpc2_same_shares_4_order2);
    assign z47_assgn47 = (temp_hpc2_v_4_order10 & a2_inp_reg);
    assign a_neg_hpc2_w_4_order10 = !a2_inp;
    assign z49_assgn49 = (a_neg_hpc2_w_4_order10_reg & rand_reg_hpc2_w_4_order10);
    assign u23 = (v23 ^ w23);
    assign z51_assgn51 = (temp_hpc2_v_4_order11 & a2_inp_reg);
    assign a_neg_hpc2_w_4_order11 = !a2_inp;
    assign z53_assgn53 = (a_neg_hpc2_w_4_order11_reg & rand_reg_hpc2_w_4_order11);
    assign u24 = (v24 ^ w24);
    assign z55_assgn55 = (temp_hpc2_v_4_order12 & a3_inp_reg);
    assign a_neg_hpc2_w_4_order12 = !a3_inp;
    assign z57_assgn57 = (a_neg_hpc2_w_4_order12_reg & rand_reg_hpc2_w_4_order12);
    assign u30 = (v30 ^ w30);
    assign z59_assgn59 = (temp_hpc2_v_4_order13 & a3_inp_reg);
    assign a_neg_hpc2_w_4_order13 = !a3_inp;
    assign z61_assgn61 = (a_neg_hpc2_w_4_order13_reg & rand_reg_hpc2_w_4_order13);
    assign u31 = (v31 ^ w31);
    assign z63_assgn63 = (temp_hpc2_v_4_order14 & a3_inp_reg);
    assign a_neg_hpc2_w_4_order14 = !a3_inp;
    assign z65_assgn65 = (a_neg_hpc2_w_4_order14_reg & rand_reg_hpc2_w_4_order14);
    assign u32 = (v32 ^ w32);
    assign z67_assgn67 = (a3_inp_reg & b_share_reg_hpc2_same_shares_4_order3);
    assign z69_assgn69 = (temp_hpc2_v_4_order15 & a3_inp_reg);
    assign a_neg_hpc2_w_4_order15 = !a3_inp;
    assign z71_assgn71 = (a_neg_hpc2_w_4_order15_reg & rand_reg_hpc2_w_4_order15);
    assign u34 = (v34 ^ w34);
    assign z73_assgn73 = (temp_hpc2_v_4_order16 & a4_inp_reg);
    assign a_neg_hpc2_w_4_order16 = !a4_inp;
    assign z75_assgn75 = (a_neg_hpc2_w_4_order16_reg & rand_reg_hpc2_w_4_order16);
    assign u40 = (v40 ^ w40);
    assign z77_assgn77 = (temp_hpc2_v_4_order17 & a4_inp_reg);
    assign a_neg_hpc2_w_4_order17 = !a4_inp;
    assign z79_assgn79 = (a_neg_hpc2_w_4_order17_reg & rand_reg_hpc2_w_4_order17);
    assign u41 = (v41 ^ w41);
    assign z81_assgn81 = (temp_hpc2_v_4_order18 & a4_inp_reg);
    assign a_neg_hpc2_w_4_order18 = !a4_inp;
    assign z83_assgn83 = (a_neg_hpc2_w_4_order18_reg & rand_reg_hpc2_w_4_order18);
    assign u42 = (v42 ^ w42);
    assign z85_assgn85 = (temp_hpc2_v_4_order19 & a4_inp_reg);
    assign a_neg_hpc2_w_4_order19 = !a4_inp;
    assign z87_assgn87 = (a_neg_hpc2_w_4_order19_reg & rand_reg_hpc2_w_4_order19);
    assign u43 = (v43 ^ w43);
    assign z89_assgn89 = (a4_inp_reg & b_share_reg_hpc2_same_shares_4_order4);
    assign t1 = (u00 ^ u01);
    assign t2 = (t1 ^ u02);
    assign t3 = (t2 ^ u03);
    assign t4 = (u10 ^ u11);
    assign t5 = (t4 ^ u12);
    assign t6 = (t5 ^ u13);
    assign t7 = (u20 ^ u21);
    assign t8 = (t7 ^ u22);
    assign t9 = (t8 ^ u23);
    assign t10 = (u30 ^ u31);
    assign t11 = (t10 ^ u32);
    assign t12 = (t11 ^ u33);
    assign t13 = (u40 ^ u41);
    assign t14 = (t13 ^ u42);
    assign t15 = (t14 ^ u43);

    always @(posedge clk) begin
        b_share_reg_hpc2_same_shares_4_order0 <= b0_inp;
        a0_inp_reg <= a0_inp;
        u00 <= z1_assgn1;
        temp_hpc2_v_4_order0 <= (b1_inp ^ r01_inp);
        v01 <= z3_assgn3;
        rand_reg_hpc2_w_4_order0 <= r01_inp;
        a_neg_hpc2_w_4_order0_reg <= a_neg_hpc2_w_4_order0;
        w01 <= z5_assgn5;
        temp_hpc2_v_4_order1 <= (b2_inp ^ r02_inp);
        v02 <= z7_assgn7;
        rand_reg_hpc2_w_4_order1 <= r02_inp;
        a_neg_hpc2_w_4_order1_reg <= a_neg_hpc2_w_4_order1;
        w02 <= z9_assgn9;
        temp_hpc2_v_4_order2 <= (b3_inp ^ r03_inp);
        v03 <= z11_assgn11;
        rand_reg_hpc2_w_4_order2 <= r03_inp;
        a_neg_hpc2_w_4_order2_reg <= a_neg_hpc2_w_4_order2;
        w03 <= z13_assgn13;
        temp_hpc2_v_4_order3 <= (b4_inp ^ r04_inp);
        v04 <= z15_assgn15;
        rand_reg_hpc2_w_4_order3 <= r04_inp;
        a_neg_hpc2_w_4_order3_reg <= a_neg_hpc2_w_4_order3;
        w04 <= z17_assgn17;
        temp_hpc2_v_4_order4 <= (b0_inp ^ r01_inp);
        a1_inp_reg <= a1_inp;
        v10 <= z19_assgn19;
        rand_reg_hpc2_w_4_order4 <= r01_inp;
        a_neg_hpc2_w_4_order4_reg <= a_neg_hpc2_w_4_order4;
        w10 <= z21_assgn21;
        b_share_reg_hpc2_same_shares_4_order1 <= b1_inp;
        u11 <= z23_assgn23;
        temp_hpc2_v_4_order5 <= (b2_inp ^ r12_inp);
        v12 <= z25_assgn25;
        rand_reg_hpc2_w_4_order5 <= r12_inp;
        a_neg_hpc2_w_4_order5_reg <= a_neg_hpc2_w_4_order5;
        w12 <= z27_assgn27;
        temp_hpc2_v_4_order6 <= (b3_inp ^ r13_inp);
        v13 <= z29_assgn29;
        rand_reg_hpc2_w_4_order6 <= r13_inp;
        a_neg_hpc2_w_4_order6_reg <= a_neg_hpc2_w_4_order6;
        w13 <= z31_assgn31;
        temp_hpc2_v_4_order7 <= (b4_inp ^ r14_inp);
        v14 <= z33_assgn33;
        rand_reg_hpc2_w_4_order7 <= r14_inp;
        a_neg_hpc2_w_4_order7_reg <= a_neg_hpc2_w_4_order7;
        w14 <= z35_assgn35;
        temp_hpc2_v_4_order8 <= (b0_inp ^ r02_inp);
        a2_inp_reg <= a2_inp;
        v20 <= z37_assgn37;
        rand_reg_hpc2_w_4_order8 <= r02_inp;
        a_neg_hpc2_w_4_order8_reg <= a_neg_hpc2_w_4_order8;
        w20 <= z39_assgn39;
        temp_hpc2_v_4_order9 <= (b1_inp ^ r12_inp);
        v21 <= z41_assgn41;
        rand_reg_hpc2_w_4_order9 <= r12_inp;
        a_neg_hpc2_w_4_order9_reg <= a_neg_hpc2_w_4_order9;
        w21 <= z43_assgn43;
        b_share_reg_hpc2_same_shares_4_order2 <= b2_inp;
        u22 <= z45_assgn45;
        temp_hpc2_v_4_order10 <= (b3_inp ^ r23_inp);
        v23 <= z47_assgn47;
        rand_reg_hpc2_w_4_order10 <= r23_inp;
        a_neg_hpc2_w_4_order10_reg <= a_neg_hpc2_w_4_order10;
        w23 <= z49_assgn49;
        temp_hpc2_v_4_order11 <= (b4_inp ^ r24_inp);
        v24 <= z51_assgn51;
        rand_reg_hpc2_w_4_order11 <= r24_inp;
        a_neg_hpc2_w_4_order11_reg <= a_neg_hpc2_w_4_order11;
        w24 <= z53_assgn53;
        temp_hpc2_v_4_order12 <= (b0_inp ^ r03_inp);
        a3_inp_reg <= a3_inp;
        v30 <= z55_assgn55;
        rand_reg_hpc2_w_4_order12 <= r03_inp;
        a_neg_hpc2_w_4_order12_reg <= a_neg_hpc2_w_4_order12;
        w30 <= z57_assgn57;
        temp_hpc2_v_4_order13 <= (b1_inp ^ r13_inp);
        v31 <= z59_assgn59;
        rand_reg_hpc2_w_4_order13 <= r13_inp;
        a_neg_hpc2_w_4_order13_reg <= a_neg_hpc2_w_4_order13;
        w31 <= z61_assgn61;
        temp_hpc2_v_4_order14 <= (b2_inp ^ r23_inp);
        v32 <= z63_assgn63;
        rand_reg_hpc2_w_4_order14 <= r23_inp;
        a_neg_hpc2_w_4_order14_reg <= a_neg_hpc2_w_4_order14;
        w32 <= z65_assgn65;
        b_share_reg_hpc2_same_shares_4_order3 <= b3_inp;
        u33 <= z67_assgn67;
        temp_hpc2_v_4_order15 <= (b4_inp ^ r34_inp);
        v34 <= z69_assgn69;
        rand_reg_hpc2_w_4_order15 <= r34_inp;
        a_neg_hpc2_w_4_order15_reg <= a_neg_hpc2_w_4_order15;
        w34 <= z71_assgn71;
        temp_hpc2_v_4_order16 <= (b0_inp ^ r04_inp);
        a4_inp_reg <= a4_inp;
        v40 <= z73_assgn73;
        rand_reg_hpc2_w_4_order16 <= r04_inp;
        a_neg_hpc2_w_4_order16_reg <= a_neg_hpc2_w_4_order16;
        w40 <= z75_assgn75;
        temp_hpc2_v_4_order17 <= (b1_inp ^ r14_inp);
        v41 <= z77_assgn77;
        rand_reg_hpc2_w_4_order17 <= r14_inp;
        a_neg_hpc2_w_4_order17_reg <= a_neg_hpc2_w_4_order17;
        w41 <= z79_assgn79;
        temp_hpc2_v_4_order18 <= (b2_inp ^ r24_inp);
        v42 <= z81_assgn81;
        rand_reg_hpc2_w_4_order18 <= r24_inp;
        a_neg_hpc2_w_4_order18_reg <= a_neg_hpc2_w_4_order18;
        w42 <= z83_assgn83;
        temp_hpc2_v_4_order19 <= (b3_inp ^ r34_inp);
        v43 <= z85_assgn85;
        rand_reg_hpc2_w_4_order19 <= r34_inp;
        a_neg_hpc2_w_4_order19_reg <= a_neg_hpc2_w_4_order19;
        w43 <= z87_assgn87;
        b_share_reg_hpc2_same_shares_4_order4 <= b4_inp;
        u44 <= z89_assgn89;
        c0 <= (t3 ^ u04);
        c1 <= (t6 ^ u14);
        c2 <= (t9 ^ u24);
        c3 <= (t12 ^ u34);
        c4 <= (t15 ^ u44);
    end

endmodule

